
`timescale 1ns/10ps
module mux32_1 (i, out, sel);
	input logic [31:0] i;
	output logic out;
	input logic [4:0] sel;
	
	logic [1:0] muxOutput;
	
	mux16_1 mux1 (.i(i[15:0]), .out(muxOutput[0]), .sel(sel[3:0]));
	mux16_1 mux2 (.i(i[31:16]), .out(muxOutput[1]), .sel(sel[3:0]));
	
	mux2_1 mux3 (.i(muxOutput), .out(out), .sel(sel[4]));
endmodule

module mux32_1_testbench ();
	logic [31:0] i;
	logic out;
	logic [4:0] sel;
	
	mux32_1 muxTest (.i, .out, .sel);
	
	initial begin
		sel=5'b01010; i = 32'b00000000000000000000010000000000; #500;
		sel=5'b00000; i = 32'b00000000000000000000000000000000; #500;   
		sel=5'b00000; i = 32'b00000001000000110111110000001001; #500;   
		sel=5'b00000; i = 32'b00000010000000110111110000001010; #500;   
		sel=5'b00000; i = 32'b00000011000000110111110000001011; #500;   
	
		sel=5'b00100; i = 32'b00001000011101111000000000000000; #500;   
		sel=5'b00100; i = 32'b00001001011101111000000000000001; #500;   
		sel=5'b00100; i = 32'b00001010011101111000000000000010; #500;   
		sel=5'b00100; i = 32'b00001011011101111000000000000100; #500;
		
		sel=5'b1011; i = 32'b01101100000111000000001001000100; #500;   
		sel=5'b1011; i = 32'b01101101001111010011111111111111; #500;   
		sel=5'b1011; i = 32'b01101110001111101110001001111000; #500;   
		sel=5'b1011; i = 32'b01101111000111110001000110000111; #500;   
		
		sel=5'b1101; i = 32'b11110001111111100000000000000111; #500;   
		sel=5'b1101; i = 32'b11110001000000000000000000000011; #500;   
		sel=5'b1101; i = 32'b11110010111100011101001100000011; #500;   
		sel=5'b1101; i = 32'b11110011110000000000110000000000; #500;  
		$finish;		
	end
endmodule
